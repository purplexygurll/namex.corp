��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  a�x�    D10      �  a�r�    D7      �  aqr    D2      �  !�+�    1      �  9�C�    0      �  	��    0      �  ����    1      �  9�C�    1      �  YQ�_    OUTPUT      �� 	 CGroupBox  Td��             �  TL�d             �  9QJ_    S3      �  9qC    1      �  !�+�    1      �  !q+    0      �  	��    1      �  	q    0      �  ����    0      �  �q�    0      �  !Q2_    S2      �  	Q_    S1      �  �Q_    S0      �  4dT�             �  d4�             �  d�             �  �d�             �  4LTd             �  L4d             �  Ld             �  �Ld             �  ����    0UNTAI MUX DENGAN 4 SELEKTOR UNTUK INPUT 2, 7, 10      �  ��i�    202031230_Rahmah Nur Fadhilah      �  1� <�     Y      �  1 )H 7    D10      �  ) � : �     D7      �  ) Q : _     D2      �  �a�o    S0      �  ya�o    S1      �  )a:o    S2      �  � a� o    S3                    ���  COR�� 	 CTerminal  h� }�               @          4�  h� }�               @          4�  �� ��               @            |� ��      5      ��    �� 	 CLogicOut4�  � �               @            � ,�      :     ��    2�4�  �� ��               @          4�  �� ��               @          4�  �� �               @            �| ��      <      ��    ��  CNAND4�  �H�I               �          4�  �X�Y              @          4�  P)Q              @            �D\     A      ��    ?�4�  �� ��                �          4�  �� ��               @          4�  � )�               @            �� �      E      ��    ?�4�  �p �q      	          �          4�  �� ��                           4�  x )y               @            �l �      I      ��    �� 	 CInverter4�  �p �q               @          4�  �p �q      	          �            �d �|      N      ��    L�4�  �� ��               @          4�  �� ��                �            �� ��      Q      ��    L�4�  �H�I     
         @          4�  �H�I               �            �<�T     T      ��    ��  CLogicIn�� 	 CLatchKey  H )X 7      W   4�  d 0y 1                            \ ,d 4     Z    ����     ��  CNAND44�  �01                          4�  �@A              @          4�  �PQ              @          4�  �`a              @          4�  DHYI     
         @            ,Dd     ]      ��8 4   [�4�  �� �                           4�  �� �               @          4�  �� �               @          4�  �� �                           4�  D� Y�               @            � D�      c      ��8 4   V�X�  @ � P �       h   4�  \ � q �                             T � \ �      j    ����     [�4�  �X Y                           4�  �h i                           4�  �x y               @          4�  �� �               @          4�  Dp Yq               @            T D�      l      ��8 4   V�X�  @ Q P _       q   4�  \ X q Y                             T T \ \      s    ����     L�4�  ��)                          4�  ����               @            ���    u      ��    L�4�  ��)                          4�  ����               @            ���    x      ��    L�4�  @A)                          4�  @�A�               @            4�L    {      ��    L�4�  � � )                          4�  � �� �               @            � �    ~      ��    V�X�  �Q�_      �   4�  �@�U                             �T�\    �    ����     V�X�  xQ�_      �   4�  �@�U                             �T�\    �    ����     V�X�  (Q8_      �   4�  @@AU                             <TD\    �    ����     V�X�  � Q� _      �   4�  � @� U                             � T� \    �    ����                   ���  CWire  �p �q      	 ��  Xp �q       ��  � 8� A       ��  � (� 9       ��  � 89      ���� 
 CCrossOver  lt      ��  ,4      ��        ��  � �         � 9       ����  >� D�       ��  �� ��       ��  �� ��         � ��       ����  ,4      ��  � ,� 4      ��  V,\4      ��  >,D4      ��  �,�4      ��  �,�4      ��  �,�4        x 0�1      ����        ��  >D      ��  V\      ��  ��      ��  ��      ��  ��        � �	      ����  � �       ��  >� D�       ��  �� ��       ��  �� ��         p � ��       ����  >� D�       ��  >D      ��  >,D4      ��  >� D�         @� Aa       ����  �� ��       ��  �� ��       ��  �� ��         �x ��        ����  �� ��       ��  ��      ��  �l�t      ��  �� ��       ��  �\�d      ��  �L�T      ��  �<�D      ��  �� ��       ��  �� ��       ��  �t �|       ��  �� ��       ��  �� ��       ��  �,�4        �h �9       ��  �� ��        ��  �� ��       ��  �� ��        ��  �� ��        ��  �� �       ��  X �      ��  X� Y       ����  lt      ��  �l�t      ��  �l�t      ��  �l�t      ��  Vl\t      ��  >lDt        � p�q      ����  � ,� 4        � � q       ��  � p� �       ����  V\      ��  Vl\t      ��  V\\d      ��  V,\4        X� Y9       ����  ��      ��  �,�4      ��  �� ��         �� �Q       ����  ��      ��  �� ��       ��  �,�4      ��  �� ��         �� �A       ��  �� �	       ��  XH�I     
 ��  �H�I      ��  �X�q       ����  �\�d      ��  �\�d      ��  �\�d      ��  V\\d        @`�a      ����  �l�t      ��  �\�d      ��  �L�T        �@��       ����  �l�t      ��  �\�d        �P��       ��  �� ��       ��  �� ��        ��  �� �       ��  hx i�        ��  (x iy       ��  @� i�       ��  @� A�        ��  (� A�       ��  @ �      ��  @ AQ       ��  (PAQ      ����  >lDt        @`A�       ��  @8Y9      ����  �� ��       ��  �� ��         �� ��       ����  �L�T      ��  �L�T        �P�Q      ����  �<�D        �@�A      ����  �� ��       ��  �� ��       ��  �� ��         X� ��       ��  �(�A       ��  @(A9       ��  @8AA       ����  �� ��       ��  �� ��         @� ��       ����  �t �|         �x �y       ��  �h �i       ����  �� ��         �� ��       ��  �8�9      ��  �(�9       ��  �8�A       ��   � 	�       ��  p X �Y                     �                            5 � 5 6 � 6 7 7 � : : < � < = � = > > A � A B � B C C E � E F � F G G � I � I J � J K K � N � N O O � Q � Q R R � T � T U U � Z Z � ] � ] ^ ^ _ _ ` � ` a a � c � c d d e e f f g g � j j � l  l m m n n o o p p � s s  u u v � v x x y � y { { | | ~ ~ �  �  � � � � � � � � � O I p N � � ~ � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � Z ] � � � � � � � � � � � � � � � � � � � � � � j c � � � � � � � � � � � � � � � � � � � � � � � � 	� � � � � � � � � J � � � � E � R Q � � � g � � � � � � � � � � � � � � � � � � �  � � � � � � � � � � � � � � � � � � � � F � a T U A B � � � � � � � � � ` � � � � � 
� v � � � � � y � < � 7 = � � 5 K � � 6 � � G �  � � C  � � | � � � � e � � � _ � � ^ � � � � f x � { � � � � o � � n � m � � d � u � > : s l             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 