��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  � �� �    C      �  � ��     V      �  )AFO    sum3      �  1ANO    sum1      �  9AVO    sum2      �  !A>O    sum0      �  �� ��     A3      �  �� ��     A2      �  �� ��     A1      �  �� ��     A0      �  �� �     F3      �  � �     F2      �  �� 	�     F1      �  �� �     F0      �  Q� ^�     M      �  � i� w    0      �  � ��    0      �  q�{�    0      �  q�{�    0      �  I�S�    0      �  ����    0      �  ����    0      �  ����    0      �  ����    0      �  ����    0      �  �i�w    0      �  �A�O    0      �  �q�    0      �  �� ��     0      �  !� +�     0      �  �� ��     0      �  '    0      �  A!K/    0      �  I!S/    0      �  9!C/    0      �  aqk    0      �  	� �     0      �  ����    0      �  ����    0      �  ��    0      �  Yg    0      �  	� �     0      �  	� �     0      �  )	3    0      �  1� ;�     0      �  � �     0      �  � �     0      �  !	+    0      �  Yqc    0      �  �Yg    0      �  y���    0      �  ����    0      �  ���    0      �  )� 3�     0      �  aikw    0      �  �i�w    0      �  ����    0      �  �I�W    0      �  ����    0      �  ����    0      �  ����    0      �  Q� [�     0      �  � �� �    1      �  9!C/    1      �  � �    1      �  ����    1      �  ����    1      �  Q�[�    1      �  ����    1      �  ����    1      �  ��    1      �  �a�o    1      �  ����    1      �  �I�W    1      �  �A�O    1      �  ��    1      �  �a�o    1      �  �I�W    1      �  �A�O    1      �  ����    1      �  ����    1      �  Q�[�    1      �  ���    1      �  ����    1      �  ���    1      �  I�S�    1      �  q�{�    1      �  q�{�    1      �  ����    1      �  ����    1      �  ���    1      �  �A�O    1      �  �q�    1      �  �� �     1      �  � #�     0      �      1      �  a �o     $UNTAI GABUNGAN FULL ADDER SUBTRACTOR      �  I� ��     202031234_M Rifqi Athallah        ����    ���  COR�� 	 CTerminal  l���     �          �          m�  l���     �          �          m�  @�U�     �          �            T�l�    n      ��    ��  CANDm�  ����     �         @          m�  ����     �          �          m�  ����     �          �            ����    s      ��    q�m�  ����     �          �          m�  ����     �                     m�  ����     �          �            ����    w      ��    �� 	 CLogicOutm�  � �� �     �          �            � x� �    |      ��    z�m�  � �� �     �         @            � �� �    ~     ��    z�m�  01-      �         @            (,8<    �     ��    ��  CXORm�  ����     �         @          m�  �x�y     �          �          m�  X�m�     �         @            lt��    �      ��    ��m�  �h�i     �          �          m�  �X�Y     �                     m�  �`�a     �          �            �T�l    �      ��    ��m�  � �� �     �         @          m�  � �� �     �          �          m�  � �� �     � 	       @            � �� �    �      ��    ��m�  � �       y                     m�  � 	�       � 	                   m�       �          �            �     �      ��    ��  CLogicIn�� 	 CLatchKey  �� ��       �   m�  �� ��      �                       �� ��     �    ����     ����  ��  �       �   m�  � 	�      �                       � �     �    ����     ��m�  (� )�       y                     m�  � �       w                     m�   !     �          �            � ,    �      ��    ��m�  �hi     �          �          m�  �XY     x         @          m�  �`�a     �         @            �T�l    �      ��    ��m�  ����     �         @          m�  �x�y     �         @          m�  h�}�     �          �            |t��    �      ��    z�m�  @A-      �          �            8,H<    �      ��    q�m�  ���     �          �          m�  ���     x         @          m�  ����     �          �            ����    �      ��    q�m�  ���     �         @          m�  ���     �         @          m�  ����     �         @            ����    �      ��    k�m�  |���     �          �          m�  |���     �         @          m�  P�e�     �         @            d�|�    �      ��    k�m�  t���     �          �          m�  t���     �         @          m�  H�]�     �         @            \�t�    �      ��    q�m�  ����     |         @          m�  ����     �         @          m�  ����     �         @            ����    �      ��    q�m�  ����     �          �          m�  ����     v         @          m�  ����     �          �            ����    �      ��    z�m�  89-      �          �            0,@<    �      ��    ��m�  ����     |         @          m�  �x�y     �         @          m�  `�u�     �          �            tt��    �      ��    ��m�  �h�i     �          �          m�  �X�Y     v         @          m�  �`�a     �         @            �T�l    �      ��    ��m�   � !�       y                     m�  � �       u                     m�       �          �            � $    �      ��    ��m�  � �       y                     m�  � 	�       t         @          m�       ~         @            �     �      ��    ��m�  �h�i     ~         @          m�  �X�Y     s         @          m�  �`�a     }          �            �T�l    �      ��    ��m�  ����     y                     m�  �x�y     }          �          m�  X�m�               �            lt��    �      ��    z�m�  01-                �            (,8<    �      ��    q�m�  ����     ~         @          m�  ����     s         @          m�  ����     z         @            ����    �      ��    q�m�  ����     y                     m�  ����     }          �          m�  ����     {          �            ����    �      ��    k�m�  l���     z         @          m�  l���     {          �          m�  @�U�     |         @            T�l�    �      ��    ����  @� P�       �   m�  0� E�      y                       D� L�     �    ����     ����  �� ��      �   m�  �� ��      x         @            �� ��     �   ����     ����   � �       �   m�  � �      w                       � �     �    ����     ����  �� ��      �   m�  �� ��      v         @            �� ��     �   ����     ����  �� �       �   m�  � �      u                       � �     �    ����     ����  ��  �      �   m�  � 	�      t         @            � �     �   ����     ����  �� ��      �   m�  �� ��      s         @            �� ��     �   ����     k�m�  � 	     _          �          m�  ��	�     ^          �          m�  ����     ]          �            ���    �      ��    q�m�  d�y�     a          �          m�  d�y�     `          �          m�  8�M�     ^          �            L�d�         ��    q�m�  dy     d          �          m�  dy	     c                     m�  8M     _          �            Ld         ��    z�m�  �1�     ]          �            ��    
     ��    z�m�  $9     e          �            $          ��    z�m�  �@�U      f          �            �T�d         ��    ��m�  �!�     a          �          m�  �!�     `          �          m�  ����     f          �            ���         ��    ��m�  d�y�     d          �          m�  d�y�     c                     m�  8�M�     `          �            L|d�         ��    ��m�  d y!     a          �          m�  dy     ]          �          m�  8M     e 	        �            Ld$         ��    ��m�  � �      g          �          m�  � �      b 	                   m�  �,�A     d          �            ��,         ��    ����  X�h�        m�  p�q	     c                       l�t�    !   ����     ����  x���      "  m�  ���     b                       ����    $   ����     ����  ��	�      %  m�  	�	�     &                       	�	�    '   ����     ����  	�(	�      (  m�  0	�1	�     $                       ,	�4	�    *   ����     ����  ��      +  m�   �!�                            �$�    -   ����     ����  (�8�      .  m�  @�A�     "                       <�D�    0   ����     ����  ���      1  m�  ��                            ��    3   ����     ����  �(�      4  m�  0�1�                            ,�4�    6   ����     ����  ����      7  m�  ����                            ����    9   ����     ����  ����      :  m�  ����                            ����    <   ����     k�m�  ����     *          �          m�  ����     +          �          m�  h�}�               �            |���    >     ��    q�m�  	�	�     (          �          m�  	�	�     '          �          m�  ����     +          �            ��	�    B     ��    q�m�  			     %          �          m�  	�	�     &                     m�  � �     *          �            ��	    F     ��    z�m�  X0YE      )          �            PD`T    J     ��    ��m�  ����     (          �          m�  ����     '          �          m�  ����     )          �            ����    L     ��    ��m�  	�	�     %          �          m�  	p	q     &                     m�  �x�y     '          �            �l	�    P     ��    ��m�  @	�A	      #          �          m�  0	�1	      $ 	                   m�  8	9	1     %          �            ,	D	    T     ��    ��m�  P�Q      !          �          m�  @�A      " 	                   m�  HI1               �            <T    X     ��    ��m�  �)�               �          m�  p)q                          m�  �x�y               �            �l�    \     ��    ��m�  ����               �          m�  ����               �          m�  ����                �            ����    `     ��    z�m�  h0iE                 �            `DpT    d     ��    q�m�  )	               �          m�  �)�                          m�  � �               �            ��    f     ��    q�m�  �)�               �          m�  �)�               �          m�  ����               �            ���    j     ��    k�m�  ����               �          m�  ����               �          m�  x���               �            ����    n     ��    k�m�  ����               �          m�  ����               �          m�  h�}�               �            |���    r     ��    q�m�  ��               �          m�  ��               �          m�  ����               �            ���    v     ��    q�m�  	               �          m�  ��                          m�  � �               �            ��    z     ��    z�m�  X0YE                �            PD`T    ~     ��    ��m�  ����               �          m�  ����               �          m�  ����               �            ����    �     ��    ��m�  ��               �          m�  pq                          m�  �x�y               �            �l�    �     ��    ��m�  @�A                �          m�  0�1       	                   m�  891               �            ,D    �     ��    ��m�   �      	          �          m�  ���       	                   m�  ��1               �            �    �     ��    ��m�  ��               �          m�  � �               �          m�  ��	      	        �            ���    �     ��    ��m�  ����               �          m�  �p�q                          m�  �x�y               �            �l��    �     ��    ��m�  l���               �          m�  l���               �          m�  @�U�     -          �            T�l�    �     ��    z�m�  0E      -          �            D T    �     ��    z�m�  ��	               �            t �    �     ��    z�m�  |���               �            l�|�    �     ��    q�m�  ��	               �          m�  ����                          m�  � �               �            ���    �     ��    q�m�  ����               �          m�  ����               �          m�  ����               �            ����    �     ��    k�m�  T�i�               �          m�  T�i�               �          m�  (�=�               �            <�T�    �     ��      ����    ���  CWire�� 
 CCrossOver  ��      ��  dl        X	�      � ��  ����      � ��  ����     � ��  ����      � ��  ����     � ��  � �� �      � ��  � �� �     � ����  .�4�        � �A�     � ��  0�Y�     � ��  ����     � ��  �x�y     � ��  �`�y      � ��  �`�a     � ��  ���     � ��  �X	Y     � ��  ��	�     � ����  dl        �hi     � ����  .�4�        � ���     � ��  ���      � ����  ����        �x��      � ��  ����      � ��  ���     � ��   ��      � ����  ����        ���     � ����  ��      ��  ��         �)�     � ��  �)     � ����  .�4�      ��  .�4�        0�1      � ��  � �� �      � ��  �� �Y      � ��  �� ��      � ����  ��        h�      � ��   !i      � ����  ����        ���     � ��   ��     � ��   ��      � ����  ����        �x��      � ����  dl         h!i     � ��   ��     x ��   �!�     � ��  �`�a     � ��  �`�y      � ��  �x�y     � ��  ���     � ��  @�i�     � ��  ����     � ��  ����      � ��  ����     � ��  ����      � ��  ����      � ��  ����     � ��  ����      � ��  ����     � ��  8�a�     � ��  ����     � ��  �x�y     � ��  �`�y      � ��  �`�a     � ��  ���     � ��  �XY     v ��  ���     v ����  dl        �hi     � ����  ����        �x��      � ��  ����      � ��  ��	�     | ����  ����        ��	�     | ��  i      � ��  i      � ��  i      ~ ����  ����        ���     y ��   ��      y ��  ���     y ��  ����      } ����  ����        �x��      } ����  dl        �hi     ~ ��  ��	�     s ��  ���     ~ ��  �`�a     } ��  �`�y      } ��  �x�y     } ��  ����     } ��  0�Y�      ��  ����     z ��  ����      z ��  ����     { ��  ����      { ��  (�)      � ����  >�D�        @�A      � ��  (�)�      � ����  >�D�        (�Q�     � ��  ��      � ����  ��      ��  dl        X�      x ����  �$�         h!�      � ����  6�<�        8�9      � ����  6�<�      ��  �$�      ��  ��        �I�     � ��  H�I�      � ��  �	�      | ����  ��      ��  dl        X�      v ����  ��        h�      � ����  .�4�        0�1       ����  .�4�      ��  ��      ��  ��        �A�     | ��  @�A�      | ��  � �       y ��  0� 1�       y ��  �� �      x ��   XY     x ����  �� �          � Y      x ����  � �         � �       w ��  (� )�       y ����  �� �       ��  � �         � )�      y ��  �� ��      v ����  �� ��         �� �Y      v ����  � �         � �       u ��   � !�       y ����  �� ��       ��  � �         (� !�      y ��  �� ��      s ��  �X	Y     s ����  �� ��         �� �Y      s ����  � �         � 	�       t ��  � �       y ����  �� ��       ��  � �          � �      y ��  � 1�      y ����  ��      ��  dl        X	�      s ����  ��        h�      ~ ����  ��      ��  ��         �1�     y ��  0� 1�      y ��  ���9      a ����  ����        ���      d ����  ����      ��  ����        ���	      c ��  �	�      ^ ��  �9�     ^ ��   	      _ ��  9     _ ��  x�y      ] ��  0�y�     ] ����  ����        x���     ] ��  ����     f ��  0�y�     ` ��   �1�     ` ��  0�1�      ` ��  0�9�     ` ��  x�     d ��  x���     c ��  x�	     c ����  ����        x���     d ����  ��$        x 	!     a ��   	9      a ����  .�4�        0�1�      ` ��  x�y�      ` ��  x���     a ��  ����      a ����  .�4�         ���     a ����  ����      ��  ����        ����     a ��  8�9     a ����  ��$      ��  ����        ���A      f ��  0�1�      ] ��  �@��      d ��  xy�      c ��  py	     c ��  	�	q      & ��  H0I�       ��  	�	�     & ��  h�i�       ����  V�\�      ��  F�L�      ��  >�D�        8�i�      ����  V�\�        X�Y1      ) ����  F�L�        H�I	       ����  >�D�      ��  >|D�        @pA�       ��  (�)q       ��   �)�      ����  f�l�        `�y�      ��  `�a�       ����  f�l�        h�i1        ����  6�<�      ��  .�4�        (�a�      ����  6�<�        8�9	       ����  .�4�      ��  .|4�        0p1�       ��  �q       ��  ��      ��  �)       ��  ��       ����  V�\�        �i�      ����  V�\�        X�Y1       ��  ����      ��  ���q       ��  ����      ��  �0��       ����  ����        ���	       ��  ����       ����        ��  ��        �1      - ��  ����      + ��  ����     + ��  ���      * ��  � �     * ��  X���     ) ��  ��	�     ' ��  ����     ' ��  �x��      ' ��  �x�y     ' ��  	9		     % ��  	p1	q     & ��  	�1	�     & ����  .	|4	�        	�9	�     % ��  8	09	�      % ��  8	�9		      % ����  ����        ����      ' ��  	�	�      ' ����  .	|4	�        0	p1	�      & ��  	�)	�     ( ��  (	�)	�      ( ����  ����        ��)	�     ( ����  ����        ��9�      ��  8�9�       ��  (�9�      ��  (�)�       ����  ����        ����       ����  >|D�        (�I�      ��  (�A�      ��  (pAq      ��  (I	      ��  �x�y      ��  �x��       ��  ����      ��  ��)�      ��  h���       ��  � �      ��  ���       ��  ����      ��  ����       ����  ����      ��  �|��        �p��       ��  ����       ��  ���       ��  � �      ��  X���      ��  ���      ��  ����      ��  �x��       ��  �x�y      ��  9	      ��  p1q      ��  �1�      ����  .|4�        �9�      ��  809�       ����  ����        ����       ��  ��       ��  �)�      ��  (�)�       ����  ����        ��)�      ��  h()      ����  ����      ��  ����        ���      ����  ����        ����      ��  ����       ��  ����      ��  ����       ����  ����        ����       ��  hi)       ����          �i      ����  �|��        ����      ��  ����      ��  �p�q      ��  ��	      ��  �x�y      ��  �x��       ��  ����      ��  ����      ��  �A�     - ����  ��        ��)�      ��  ����      ��  ���       ��  h �      ��  h�i       ��  h���      ��  h�i�         ����    �  ����      ����    n n �o o �p �p s s �t t �u �u w w �x x �y �y | | �~ ~ � � �� � � �� � �� �� � � �� � �� �� � � �� � �� ~ � � :� � � � � � � � �� � � � B� � @� � � �� � �� � =� �� � � �� � �� �� � � � � �� � �� �� � � �� � �� �� � � �� � �� � � � �� � �� ,� � �  � � �� �� � � �� � �� �� � &� � � � � �� �� � � �� � �� �� � K� � I� � � � U� � S� � � � � � � P� � � � � � � � � 3� � � � � � � � � 	� � 
� � � � � � � 9� � ;� � � <� � @� � F� � I� � S� � O� � k� � i o ��jvxl

���sqywu{m  $�!!�$$''�**U--�00Y33�66�99�<<�>>�??�@�@BB�CC�D�DFF�GG�H�HJ�JLL�MM�N�NPP�QQ�R�RT  TU*UVV�X  XY0YZZ�\\�]]�^�^``�aa�b�bd�dff�gg�h�hjj�kk�l�lnn�oo�p�prr�ss�t�tvvwwx�xzz�{{�|�|~�~������������������  ��6�����  ��9��������!�����������
������������������"������$���#��%���������o �u n ��y �� �����p �� ��� ����� w ���x ���� ���� ��������t s ������ ������������� | ��� � ����� ���� (�  �� �����#� $� !� $�� ��� ���� �� � ��� �� �� �� � ��� &� ��� ����� � 1G.� .�0� 1����� � -�� -� �� �� � _	� � \� ]� Z� ]� � 
3� � � � � ��� �� ��!+!�=�$*��&)�� ('(%(" ,(� 5 .8.���17�36� 54525/95� C� Yb� >>!>D<� @E� � L� C?CA:B� GGMF� IN� � V� LHLJCK� QQZQWO� SX� � Y� VRVTLUV;ZaZP]`_^_[b� _��d��vf�fzwxj� i� lko�mo�n �~�~ustd�ffyhd{�}{�~�trr������g�e�c}c�|�pq
ny�!��QZ�'��@�����������J�����������]-����p�����d�����������������3������t���~<����x��	�� ����?�D>��H�N��M����RF���G���P�V��������C����B�����L���`���j��k������\�g���f��^��a����b�hn��l�o���sr��|���������z���{�����������wv �����
�
������������������� ��!�#��"%�$� �          �$s�        @     +        @            @    "V  (      H	x                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 