��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  9)P7    A10      �  9	J    A7      �  9�J�    A2      �� 	 CGroupBox  ,�d@             �  ����             �  ����             �  ���             �  �,�             �  ���@             �  ���@             �  ��@             �  �,@             �  ����    F0      �  ����    F1      �  ��	�    F2      �  ����    0      �  �	�    0      �  ����    0      �  �	�    1      �  ���    0      �  �	    1      �  ��    1      �  �!�    F3      �  ,�d�             �  1�`�    OUTPUT      �  	    1      �  �)�7    1      �  �)�7    0      �  )7    0      �  �)7    1      �  YQ �_     UNTAI MUX 4 SELEKTOR  2,7,10      �  	Y g    A10      �  	�     A7      �  i�y�    F3      �  ����    F2      �  ��    F1      �  I�Y�    F0      �  i� t�     Y      �  	� �     A2      �  �� N�     202031234_M Rifqi Athallah                    ���  CLogicIn�� 	 CLatchKey   Y0g      3   �� 	 CTerminal  <`Qa                            4\<d     7    ����     2�4�   � 0      8   6�  < Q                            4� <     :    ����     2�4�  hqx      ;   6�  �`�u       	                     |t�|    =    ����     2�4�  �q�      >   6�  �`�u       	                     �t�|    @    ����     2�4�   q      A   6�  `u       	                     t|    C    ����     2�4�  HqX      D   6�  ``au       	                     \td|    F    ����     �� 	 CInverter6�  La                          6�   5               @            4$L    I      ��    G�6�  `Laa                          6�  ` a5               @            T4lL    L      ��    ��  CNAND46�  �� ��               @          6�  �� ��                           6�  �� ��               @          6�  �� ��               @          6�  �� 	�               @            �� ��      P      ��8 4   G�6�  � �       	       @          6�  4� I�                �            � 4�      V      ��    ��  CAND6�  H� ]�       	        �          6�  H� ]�                           6�  t� ��      	          �            \� t�      Z      ��    N�6�  �`�a                          6�  �p�q              @          6�  ����              @          6�  ����              @          6�  �x	y              @            �\��     ^      ��8 4   G�6�  xy      	       @          6�  4xIy               �            l4�     d      ��    X�6�  Hx]y      	        �          6�  H�]�              @          6�  t���               �            \tt�     g      ��    N�6�  � �                          6�  ��              @          6�  � �!              @          6�  �0�1                          6�  �	              @            �� �4     k      ��8 4   G�6�        	       @          6�  4I               �            4$     q      ��    X�6�  H]      	        �          6�  H(])              @          6�  t �!     
          �            \t,     t      ��    ��  COR6�  �� ��      	          �          6�  �� ��      
          �          6�  �� ��                �            �� ��      y      ��    w�6�  �� �                �          6�  �� �                �          6�  � 1�                �            � �      }      ��    �� 	 CLogicOut6�  @� U�                �            T� d�      �      ��    2�4�   � 0�      �   6�  <� Q�               @            4� <�      �   ����     G�6�  �L�a                          6�  � �5               @            t4�L    �      ��    G�6�  �L�a                          6�  � �5               @            �4�L    �      ��                  ���  CWire  �� ��       ��  �� ��       ��  ����      ��  �� ��      
 ��  �� �!      
 ��  �� ��      	 ��  �� ��       ��  0� A�       ��  P� ��       ��  x� ��       ��  ``ya      ���� 
 CCrossOver  v� |�         � ��       ����  � �       ��  v� |�         �� ��       ��  �� I�       ��  �� ��        ����  �� ��       ��  � �       ��  v� |�         �� ��       ����  �� �      ��  �� �      ��  �       ��  v� |        P �      ��  �`�a      ����  v|        `�      ����  ^d$      ��  v|$         �!      ����  �       ��  � �       ��  � �         � !       ����  ,4      ��  ^,d4      ��  v,|4        �0�1      ��  �`�a      ��   (I)      ��   (A       ����  ~\�d      ��  �\�d      ��  ^\dd      ��  �\�d      ��  �\�d      ��  \d      ��  v\|d        P`�a      ����  �<�D      ��  �<�D      ��  �<�D      ��  <D      ��  ^<dD      ��  v<|D        �@A      ����  vl|t        `p�q      ����  ^\dd      ��  ^d$      ��  ^,d4      ��  ^<dD        `aq       ����  ^|d�      ��  v||�        ���      ����  \d      ��  ,4      ��  <D         �       ����  ����      ��  ��      ��  ^�d�      ��  v�|�        ����      ����  �� �      ��  �\�d      ��  �� ��       ��  �<�D        �� ��       ��  ��I�      ����  v�|�      ��  v�|�      ��  v||�      ��  vl|t      ��  v<|D      ��  v,|4      ��  v|$      ��  v|      ��  v� |�       ��  v� |�       ��  v� |�       ��  v\|d      ��  v� |        x� ya       ����  ^�d�      ��  ^�d�      ��  ^|d�        `pa!       ����  ��      ��  ��        �!       ����  ����      ��  ����      ��  �<�D      ��  �\�d        �0�a       ����  ����        ���!       ����  ����      ��  �<�D      ��  �\�d      ��  �� �        �� �a       ��  ����       ����  ����      ��  ����      ��  ����      ��  ��      ��  ^�d�      ��  v�|�        ����      ����  ~\�d        �@��       ��  ���!                     �                            7 7 � : : � = � = @ � @ C I C F � F I I C J � J L L F M � M P � P Q � Q R � R S � S T T V V T V W W Z Z W Z [ � [ \ \ � ^ � ^ _ � _ ` � ` a � a b b d d b d e e g g e g h � h i i � k � k l � l m � m n � n o o q q o q r r t t r t u � u v v � y � y z � z { { � } � } ~ � ~   � � � � � � � � � = � � � � @ � � � � ~ � � i � � z � v \ y { }  � � P � Q L � � � � R � � � � � S � [ � � � � � � � � � � � � � � � � � : k � � � � � l � � � � � m � � � � � � � � � � � � � � � n � � � u � � � � � � � � � � � � � � 7 ^ � � � � � � � � � � � � � � � _ � � � � � � � � � � � � � � � ` � � � � � � � � � � � � � � � � � a � � � � � � � � � � h � � � � � � � � � � � � � � � � � � � � � � � � � � � � 
� � � � � M � 	� � � J � � � � � � � � � � � � � � � � � � � � � �  � � � � � � � �             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 